library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

-- THIS IS TO CHOOSE THE TYPE OF IMMEDIATE EXTENSION -- ZERO OR SIGNED
-- ExtOp is the selection bit


ENTITY SEFA_IMMEDIATE_EXTENDED_MUX IS
PORT(
		SEFA_ZERO_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGN_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_ExtOp : IN STD_LOGIC;
		SEFA_EXTENDED_IMM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_IMMEDIATE_EXTENDED_MUX;

ARCHITECTURE ARCH OF SEFA_IMMEDIATE_EXTENDED_MUX IS
	
BEGIN


	SEFA_EXTENDED_IMM <= SEFA_SIGN_EXTENDED_IMM WHEN SEFA_ExtOp = '1' 
							ELSE SEFA_ZERO_EXTENDED_IMM;

END ARCH;
