LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

-- THE PURPOSE OF THIS VALUE IS TO SAVE THE CURRENT PC VALUE. 
-- WILL ADD MORE DETAILS LATER AS IT CONNECTS. 

ENTITY SEFA_STORE_PC_VALUE IS
PORT(
	SEFA_CLOCK: IN STD_LOGIC;
	SEFA_PC_INPUT: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_PC_OUTPUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_STORE_PC_VALUE;

ARCHITECTURE ARCH OF SEFA_STORE_PC_VALUE IS
	SIGNAL SEFA_PC_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	BEGIN
		PROCESS(SEFA_CLOCK)
		BEGIN
			IF(RISING_EDGE(SEFA_CLOCK)) THEN
					SEFA_PC_OUT <= SEFA_PC_INPUT; --UPDATE CURRENT PC VALUE. 
			END IF;
		END PROCESS;
		SEFA_PC_OUTPUT <= SEFA_PC_OUT;
END ARCH;
	