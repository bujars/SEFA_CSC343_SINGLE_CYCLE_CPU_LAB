LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE SEFA_SINGLE_CYCLE_CPU_PACKAGE IS

COMPONENT SEFA_ALU IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
--	SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
--	SEFA_FUNCT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_ALUctr : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ALU_OUTPUT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_HI : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_LO : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
	
	-- NOTE IM NOT SURE HOW WE ARE GOING TO DO OUTPUT FOR MUL/DIV WHICH IS 64 BITS.......FOR NOW IGNORING.
);
END COMPONENT SEFA_ALU;

COMPONENT SEFA_ALU_MUX IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
--	SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
--	SEFA_FUNCT: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_ALUctr : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	SEFA_ADD : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_SUB : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ADDU : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ADDI : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ADDIU : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_SUBU : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_AND : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_OR : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_NOR : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ANDI : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ORI : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_MULT : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
	SEFA_DIVIDE_QUOTIENT : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_DIVIDE_REMAINDER : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ALU_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
	-- NOTE IM NOT SURE HOW WE ARE GOING TO DO OUTPUT FOR MUL/DIV WHICH IS 64 BITS.......FOR NOW IGNORING.
);
END COMPONENT SEFA_ALU_MUX;

COMPONENT SEFA_SIGNED_LPM_ADD_SUB IS
	PORT
	(
		SEFA_add_sub		: IN STD_LOGIC ;
		SEFA_dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_overflow		: OUT STD_LOGIC ;
		SEFA_result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_SIGNED_LPM_ADD_SUB;

COMPONENT SEFA_UNSIGNED_LPM_ADD_SUB IS
	PORT
	(
		SEFA_add_sub		: IN STD_LOGIC ;
		SEFA_dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_UNSIGNED_LPM_ADD_SUB;

COMPONENT SEFA_AND_COMPONENT IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_AND_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
);
END COMPONENT SEFA_AND_COMPONENT;

COMPONENT SEFA_OR_COMPONENT IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_OR_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
);
END COMPONENT SEFA_OR_COMPONENT;

COMPONENT SEFA_NOR_COMPONENT IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_NOR_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
);
END COMPONENT SEFA_NOR_COMPONENT;

COMPONENT SEFA_LPM_MULT IS
	PORT
	(
		SEFA_dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
END COMPONENT SEFA_LPM_MULT;

COMPONENT SEFA_LPM_DIVIDE IS
	PORT
	(
		SEFA_denom		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_numer		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_quotient		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_remain		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_LPM_DIVIDE;


COMPONENT SEFA_Register_N_VHDL is 
	generic (SEFA_N: integer := 32); -- The genetics feature permits us to change the side of this register desin easily. Its a const variable
	port (
		SEFA_clk: in std_logic; -- clock
		SEFA_wren: in std_logic; -- write enable (if it is 0, the stored data will not change)
		SEFA_rden: in std_logic; -- read enable (only when it is 1, the stored data will be displayed to output)
		SEFA_chen: in std_logic; --  chip enable (if it is 0, the output will be undefined)
		SEFA_data: in std_logic_vector (SEFA_N-1 downto 0); -- data input
		SEFA_q: out std_logic_vector(SEFA_N-1 downto 0) -- output. This is essentially just a display
		);
end COMPONENT SEFA_Register_N_VHDL;


COMPONENT SEFA_IR_REGISTER IS
	generic (SEFA_N: integer := 32);
	port(
	SEFA_clk: in std_logic; -- clock
		SEFA_wren: in std_logic; -- write enable (if it is 0, the stored data will not change)
		SEFA_rden: in std_logic; -- read enable (only when it is 1, the stored data will be displayed to output)
		SEFA_chen: in std_logic; --  chip enable (if it is 0, the output will be undefined)
		SEFA_data: in std_logic_vector (SEFA_N-1 downto 0); -- data input
		SEFA_IR: out std_logic_vector(SEFA_N-1 downto 0)
		);
end COMPONENT SEFA_IR_REGISTER;

COMPONENT SEFA_PC_REGISTER IS
	generic (SEFA_N: integer := 32);
	port(
	SEFA_clk: in std_logic; -- clock
		SEFA_wren: in std_logic; -- write enable (if it is 0, the stored data will not change)
		SEFA_rden: in std_logic; -- read enable (only when it is 1, the stored data will be displayed to output)
		SEFA_chen: in std_logic; --  chip enable (if it is 0, the output will be undefined)
		SEFA_data: in std_logic_vector (SEFA_N-1 downto 0); -- data input
		SEFA_PC: out std_logic_vector(SEFA_N-1 downto 0)
		);
end COMPONENT SEFA_PC_REGISTER;

COMPONENT SEFA_PC_PLUS_4 IS
	PORT(
		SEFA_PC_OLD : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_PC_NEW : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT SEFA_PC_PLUS_4;

COMPONENT SEFA_PC_PLUS_IMMEDIATE_PLUS_4 IS
	PORT(
		SEFA_PC_PLUS_4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGN_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_PC_NEW : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT SEFA_PC_PLUS_IMMEDIATE_PLUS_4;


COMPONENT SEFA_SIGN_EXTEND_IMM_16_TO_32 IS
PORT (
		SEFA_IMM16 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		SEFA_IMM32 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_SIGN_EXTEND_IMM_16_TO_32;

COMPONENT SEFA_ZERO_EXTEND_IMM_16_TO_32 IS
PORT (
		SEFA_IMM16 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		SEFA_IMM32 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_ZERO_EXTEND_IMM_16_TO_32;

COMPONENT SEFA_SIGN_EXTEND_IMM_26_TO_32 IS
PORT (
		SEFA_IMM26 : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
		SEFA_IMM32 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_SIGN_EXTEND_IMM_26_TO_32;

COMPONENT SEFA_BRANCHING_MUX IS
	PORT(
		SEFA_PCSrc : IN STD_LOGIC;
		SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		SEFA_PC_Plus_4 : IN STD_LOGIC_VECTOR(31 DOWNTo 0);
		SEFA_PC_IMM_Plus_4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_PC_SELECTOR : IN STD_LOGIC; 
		SEFA_PC_NEW : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT SEFA_BRANCHING_MUX;

COMPONENT SEFA_BRANCHING_SIGNED_EXTENDED IS
PORT(
		SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		SEFA_SIGNED_16_to_32_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGNED_26_to_32_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGNED_32_EXTENDED_IMM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_BRANCHING_SIGNED_EXTENDED;

COMPONENT SEFA_SELECT_SECOND_ALU_INPUT IS
PORT(
		SEFA_BUSB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_ALUsrc : IN STD_LOGIC;
		SEFA_INPUT_B : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_SELECT_SECOND_ALU_INPUT;

COMPONENT SEFA_IMMEDIATE_EXTENDED_MUX IS
PORT(
		SEFA_ZERO_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGN_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_ExtOp : IN STD_LOGIC;
		SEFA_EXTENDED_IMM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_IMMEDIATE_EXTENDED_MUX;

COMPONENT SEFA_IMMEDIATE_EXTENDER IS
PORT(
		SEFA_IMM16 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		SEFA_ExtOp : IN STD_LOGIC;
		SEFA_EXTENDED_IMM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_IMMEDIATE_EXTENDER;


COMPONENT SEFA_CPU_CONTROL_SIGNALS IS
PORT(
	SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0); -- NOTE I MIGHT BE ABLE TO SIMPLIFY THIS TO JUST OPCODE OR FUNCT AS WE DON'T HAVE MIXED VALUES AS OF NOW...
	SEFA_FUNCT: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_ALUctr : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	SEFA_ExtOp : OUT STD_LOGIC;
	SEFA_ALUSrc : OUT STD_LOGIC;
	SEFA_MemWr : OUT STD_LOGIC;
	SEFA_MemtoReg : OUT STD_LOGIC;
	SEFA_PCSrc : OUT STD_LOGIC;
	SEFA_RegDst : OUT STD_LOGIC;
	SEFA_RegWr : OUT STD_LOGIC

);
END COMPONENT SEFA_CPU_CONTROL_SIGNALS;


COMPONENT SEFA_RAM3PORT IS
PORT
(
	SEFA_clock : IN STD_LOGIC;
	SEFA_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	SEFA_rdaddress_a : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	SEFA_rdaddress_b : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	SEFA_wraddress : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	SEFA_wren : IN STD_LOGIC := '1';
	SEFA_qa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
	SEFA_qb : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
);

END COMPONENT SEFA_RAM3PORT;

COMPONENT SEFA_DATA_MEMORY_RAM_1_PORT IS
	PORT
	(
		SEFA_address		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		SEFA_clock		: IN STD_LOGIC  := '1';
		SEFA_data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_wren		: IN STD_LOGIC ;
		SEFA_q		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_DATA_MEMORY_RAM_1_PORT;


COMPONENT SEFA_INSTRUCTION_MEMORY_RAM_1_PORT IS
	PORT
	(
		SEFA_address		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		SEFA_clock		: IN STD_LOGIC  := '1';
		SEFA_data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_wren		: IN STD_LOGIC ;
		SEFA_q		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_INSTRUCTION_MEMORY_RAM_1_PORT;

COMPONENT SEFA_SELECT_MEM_TO_REG IS
PORT(
		SEFA_ALU_OUTPUT: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_DATA_MEM_OUTPUT : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_MemtoReg : IN STD_LOGIC;
		SEFA_MEM_TO_REG_OUTPUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_SELECT_MEM_TO_REG;

COMPONENT SEFA_SELECT_REGISTER_FILE_INPUT IS
PORT(
		SEFA_RT: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		SEFA_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		SEFA_RegDst : IN STD_LOGIC;
		SEFA_REGISTER_FILE_SELECTED_INPUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
);
END COMPONENT SEFA_SELECT_REGISTER_FILE_INPUT;


--COMPONENT SEFA_IR_DRIVER IS 
--GENERIC(SEFA_N : INTEGER := 32);
--PORT(
--	SEFA_CLOCK : IN STD_LOGIC; --- NEED TO ADD CLOCK AS INPUT.
--	SEFA_IR_INPUT : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
--	-- SEFA_SOME_UNKNOWN_OUTPUT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0) -- ONLY USED FOR TESTING PURPOSES.
--);
--END COMPONENT SEFA_IR_DRIVER;


COMPONENT SEFA_IR_DRIVER IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_CLOCK : IN STD_LOGIC; --- NEED TO ADD CLOCK AS INPUT. 
	--SEFA_IR_INPUT : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	-- SEFA_SOME_UNKNOWN_OUTPUT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0) -- THIS WAS ONLY USED FOR TESTING PURPOSES.
	
	SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0); -- ALL INSTRUCTION
	SEFA_RS : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SEFA_RT : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SEFA_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SEFA_SHAMT : IN STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SEFA_FUNCT :  IN STD_LOGIC_VECTOR(5 DOWNTO 0); -- R INSTRUCTION
	SEFA_IMM16 :  IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- I INSTRUCTION
	SEFA_IMM26 : IN STD_LOGIC_VECTOR(25 DOWNTO 0); -- J INSTRUCTION
	SEFA_ALUctr : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	SEFA_ExtOp : IN STD_LOGIC;
	SEFA_ALUSrc : IN STD_LOGIC;
	SEFA_MemWr : IN STD_LOGIC;
	SEFA_MemtoReg : IN STD_LOGIC;
	SEFA_PCSrc : IN STD_LOGIC;
	SEFA_RegDst : IN STD_LOGIC;
	SEFA_RegWr : IN STD_LOGIC
	
	
	
	
);
END COMPONENT SEFA_IR_DRIVER;

COMPONENT SEFA_NON_LPM_REGISTER_FILE IS
PORT(
	SEFA_clock: IN STD_LOGIC;
	SEFA_data: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_wraddress: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	SEFA_rdaddress_a: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	SEFA_rdaddress_b: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	SEFA_wren: IN STD_LOGIC;
	SEFA_qa: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_qb: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_NON_LPM_REGISTER_FILE;


COMPONENT SEFA_NON_LPM_DATA_MEMORY IS
PORT(
	SEFA_clock: IN STD_LOGIC;
	SEFA_data: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_address: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	SEFA_wren: IN STD_LOGIC;
	SEFA_q: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_NON_LPM_DATA_MEMORY;

COMPONENT SEFA_NON_LPM_INSTRUCTION_MEMORY IS
PORT(
	SEFA_clock: IN STD_LOGIC;
	SEFA_data: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_address: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	SEFA_wren: IN STD_LOGIC;
	SEFA_q: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_NON_LPM_INSTRUCTION_MEMORY;



COMPONENT SEFA_STORE_PC_VALUE IS
PORT(
	SEFA_CLOCK: IN STD_LOGIC;
	SEFA_PC_INPUT: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_PC_OUTPUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_STORE_PC_VALUE;

COMPONENT SEFA_Comparator_N IS
	GENERIC(SEFA_N : INTEGER := 32);
	PORT(
			SEFA_IN0, SEFA_IN1 : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
			SEFA_OUT : OUT STD_LOGIC
	);
end COMPONENT SEFA_Comparator_N;


COMPONENT SEFA_NAL IS
PORT(
		SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0); -- KEEPING BECAUSE HASSLE TO CHANGE. 
		SEFA_PCSrc : IN STD_LOGIC;
		SEFA_PC_COND : IN STD_LOGIC;
		SEFA_PC_OLD : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_IMM16 : IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- NOTE THIS IS 16 BITS AND WE NEED TO SIGN EXTEND! 
		SEFA_IMM26 : IN STD_LOGIC_VECTOR(25 DOWNTO 0); -- NOTE THIS IS 26 BITS AND WE NEED TO SIGN EXTEND! 
		SEFA_UPDATED_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END COMPONENT SEFA_NAL;

COMPONENT SEFA_MAIN IS PORT(
	SEFA_CLOCK : IN STD_LOGIC
);
END COMPONENT SEFA_MAIN;

COMPONENT SEFA_HI_REGISTER IS
	generic (SEFA_N: integer := 32);
	port(
	SEFA_clk: in std_logic; -- clock
		SEFA_wren: in std_logic; -- write enable (if it is 0, the stored data will not change)
		SEFA_rden: in std_logic; -- read enable (only when it is 1, the stored data will be displayed to output)
		SEFA_chen: in std_logic; --  chip enable (if it is 0, the output will be undefined)
		SEFA_data: in std_logic_vector (SEFA_N-1 downto 0); -- data input
		SEFA_HI: out std_logic_vector(SEFA_N-1 downto 0)
		);
end COMPONENT SEFA_HI_REGISTER;

COMPONENT SEFA_LO_REGISTER IS
	generic (SEFA_N: integer := 32);
	port(
	SEFA_clk: in std_logic; -- clock
		SEFA_wren: in std_logic; -- write enable (if it is 0, the stored data will not change)
		SEFA_rden: in std_logic; -- read enable (only when it is 1, the stored data will be displayed to output)
		SEFA_chen: in std_logic; --  chip enable (if it is 0, the output will be undefined)
		SEFA_data: in std_logic_vector (SEFA_N-1 downto 0); -- data input
		SEFA_LO: out std_logic_vector(SEFA_N-1 downto 0)
		);
end COMPONENT SEFA_LO_REGISTER;


END SEFA_SINGLE_CYCLE_CPU_PACKAGE;