library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

-- THIS IS TO CHOOSE THE APPROPRIATE IMMEDIATE NUMBER OF BITS TO EXTEND (I VS J)
-- NOTE THE OPCODE 2HEX IS FOR JUMP INSTRUCTION IN THE GREEN PAGES https://courses.cs.washington.edu/courses/cse378/09au/MIPS_Green_Sheet.pdf


ENTITY SEFA_BRANCHING_SIGNED_EXTENDED IS
PORT(
		SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		SEFA_SIGNED_16_to_32_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGNED_26_to_32_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_SIGNED_32_EXTENDED_IMM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_BRANCHING_SIGNED_EXTENDED;

ARCHITECTURE arch OF SEFA_BRANCHING_SIGNED_EXTENDED IS
	
BEGIN


	SEFA_SIGNED_32_EXTENDED_IMM <= SEFA_SIGNED_26_to_32_EXTENDED_IMM WHEN SEFA_OPCODE = "000010" 
							ELSE SEFA_SIGNED_16_to_32_EXTENDED_IMM;

END arch;

