LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.ALL;

-- SWITCHING OVER TO HARDCODED BECAUSE LPM IS GIVING ME ISSUES.


ENTITY SEFA_NON_LPM_REGISTER_FILE IS
PORT(
	SEFA_clock: IN STD_LOGIC;
	SEFA_data: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_wraddress: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	SEFA_rdaddress_a: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	SEFA_rdaddress_b: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	SEFA_wren: IN STD_LOGIC;
	SEFA_qa: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_qb: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_NON_LPM_REGISTER_FILE;


ARCHITECTURE ARCH OF SEFA_NON_LPM_REGISTER_FILE IS
	TYPE SEFA_REGISTERS IS ARRAY(0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_MEM: SEFA_REGISTERS := (
	 OTHERS => X"00000000"
	);	
BEGIN
	PROCESS(SEFA_clock)
	 BEGIN
		IF (SEFA_clock'EVENT AND SEFA_clock = '1') THEN
			IF(SEFA_wren = '1') THEN
				SEFA_MEM(TO_INTEGER(UNSIGNED(SEFA_wraddress))) <= SEFA_data;
		END IF;
	END IF;
	END PROCESS;
	SEFA_qa <= SEFA_MEM(TO_INTEGER(UNSIGNED(SEFA_rdaddress_a)));
	SEFA_qb <= SEFA_MEM(TO_INTEGER(UNSIGNED(SEFA_rdaddress_b)));
END ARCH;