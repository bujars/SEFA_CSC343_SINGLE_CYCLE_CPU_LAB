LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

ENTITY SEFA_MAIN IS PORT(
	SEFA_CLOCK : IN STD_LOGIC
);
END SEFA_MAIN;


ARCHITECTURE SYN OF SEFA_MAIN IS 

		
		SIGNAL SEFA_PC : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0'); 
		-- THIS IS THE PROGRAM COUNTER VALUE.
		-- WE DEFAULT IT AT 0, AND WILL START AT 0. 

		SIGNAL SEFA_PC_NEXT: STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		
		--INSTRUCTION
		SIGNAL SEFA_INSTRUCTION : STD_LOGIC_VECTOR(31 DOWNTO 0);
		SIGNAL SEFA_IR_INSTRUCTION : STD_LOGIC_VECTOR(31 DOWNTO 0);
		
		
		SIGNAL SEFA_INSTRUCTION_ADDRESS : STD_LOGIC_VECTOR(4 DOWNTO 0);
		
		
			-- JUST FOR CLEANESS, I MIGHT MOVE THIS TO ITS OWN FILE TO SPLIT COMPONENTS. 
	SIGNAL SEFA_OPCODE : STD_LOGIC_VECTOR(5 DOWNTO 0); -- ALL INSTRUCTION
	SIGNAL SEFA_RS : STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SIGNAL SEFA_RT : STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SIGNAL SEFA_RD : STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SIGNAL SEFA_SHAMT : STD_LOGIC_VECTOR(4 DOWNTO 0); -- R INSTRUCTION
	SIGNAL SEFA_FUNCT : STD_LOGIC_VECTOR(5 DOWNTO 0); -- R INSTRUCTION
	SIGNAL SEFA_IMM16 : STD_LOGIC_VECTOR(15 DOWNTO 0); -- I INSTRUCTION
	SIGNAL SEFA_IMM26 : STD_LOGIC_VECTOR(25 DOWNTO 0); -- J INSTRUCTION
	SIGNAL SEFA_ALUctr : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL SEFA_ExtOp : STD_LOGIC;
	SIGNAL SEFA_ALUSrc : STD_LOGIC;
	SIGNAL SEFA_MemWr : STD_LOGIC;
	SIGNAL SEFA_MemtoReg : STD_LOGIC;
	SIGNAL SEFA_PCSrc : STD_LOGIC;
	SIGNAL SEFA_RegDst : STD_LOGIC;
	SIGNAL SEFA_RegWr : STD_LOGIC;
	
	-- comparator result
	SIGNAL SEFA_PC_COND : STD_LOGIC; 
	
	
	SIGNAL SEFA_REGISTER_FILE_SELECTED_INPUT : STD_LOGIC_VECTOR(4 DOWNTO 0);
	
	
	
	SIGNAL SEFA_BUS_A : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_BUS_B : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_BUS_W : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	
	SIGNAL SEFA_EXTENDED_IMM : STD_LOGIC_VECTOR(31 DOWNTO 0);

	
	SIGNAL SEFA_INPUT_B : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	
	
	--- NOTE THIS WILL CHANGE ONCE WE INCORPERATE MULTIPLY AND DIVIDE!
	SIGNAL SEFA_ALU_OUTPUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL SEFA_HI : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_LO : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL SEFA_HI_REGISTER_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SEFA_LO_REGISTER_VALUE : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	
	
	SIGNAL SEFA_DATA_MEM_OUTPUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
		
		
	
	

BEGIN
	

	GET_CURRENT_PC: SEFA_STORE_PC_VALUE PORT MAP(
			SEFA_CLOCK => SEFA_CLOCK,  
			SEFA_PC_INPUT => SEFA_PC_NEXT,
			SEFA_PC_OUTPUT => SEFA_PC
	); 
		
	
	SEFA_INSTRUCTION_ADDRESS <= SEFA_PC(6 DOWNTO 2);
	
	
	GET_INSTRUCTION_MEMORY: SEFA_NON_LPM_INSTRUCTION_MEMORY PORT MAP(
			SEFA_clock => SEFA_CLOCK,
			SEFA_data => X"00000000", -- WE ARENT STORING ANYTHING
			SEFA_address => SEFA_INSTRUCTION_ADDRESS,
			SEFA_wren => '0', -- WE ARENT WRITING ANYTHING. 
			SEFA_q => SEFA_INSTRUCTION	
	);
	
	
	PUT_INSTRUCTION_IN_IR: SEFA_IR_REGISTER PORT MAP (
		SEFA_clk => SEFA_CLOCK,
		SEFA_wren => '1',
		SEFA_rden => '1',
		SEFA_chen => '1',
		SEFA_data => SEFA_INSTRUCTION, 
		SEFA_IR => SEFA_IR_INSTRUCTION
		);
		
		
		
	-- possibly put all of this in a seperate file like the last lab. 
	SEFA_OPCODE <= SEFA_IR_INSTRUCTION(31 DOWNTO 26);
	SEFA_RS <= SEFA_IR_INSTRUCTION(25 DOWNTO 21);
	SEFA_RT <= SEFA_IR_INSTRUCTION(20 DOWNTO 16);
	SEFA_RD <= SEFA_IR_INSTRUCTION(15 DOWNTO 11);
	SEFA_SHAMT <= SEFA_IR_INSTRUCTION(10 DOWNTO 6);
	SEFA_FUNCT <= SEFA_IR_INSTRUCTION(5 DOWNTO 0);
	SEFA_IMM16 <= SEFA_IR_INSTRUCTION(15 DOWNTO 0);
	SEFA_IMM26 <= SEFA_IR_INSTRUCTION(25 DOWNTO 0);
	
	
	SET_CONTROL_SIGNALS: SEFA_CPU_CONTROL_SIGNALS PORT MAP (
											SEFA_OPCODE => SEFA_OPCODE,
											SEFA_FUNCT => SEFA_FUNCT,
											SEFA_ExtOp => SEFA_ExtOp,
											SEFA_ALUctr => SEFA_ALUctr,
											SEFA_ALUSrc => SEFA_ALUSrc,
											SEFA_MemWr => SEFA_MemWr,
											SEFA_MemtoReg => SEFA_MemtoReg,
											SEFA_PCSrc => SEFA_PCSrc,
											SEFA_RegDst => SEFA_RegDst,
											SEFA_RegWr => SEFA_RegWr
	);
		
		
		
		
--		
--		
--		MOVING ALL OF THIS INTO ONE FILE BECAUSE OF BEQ AND BNE. 
-- 	ITS REQUIRING THE VALUES OF BUS A (RS) AND BUS B (RT) WHICH WE NEED FROM IR_DRIVER. 
--		
--		
--	IR_DRIVER : SEFA_IR_DRIVER PORT MAP (
--			SEFA_CLOCK => SEFA_CLOCK, 
--			SEFA_IR_INPUT => SEFA_IR_INSTRUCTION
--			SEFA_OPCODE => SEFA_OPCODE,
--			SEFA_RS => SEFA_RS, 
--			SEFA_RT => SEFA_RT,
--			SEFA_RD => SEFA_RD, 
--			SEFA_SHAMT => SEFA_SHAMT, 
--			SEFA_FUNCT => SEFA_FUNCT, 
--			SEFA_IMM16 => SEFA_IMM16, 
--			SEFA_IMM26 => SEFA_IMM26, 
--			SEFA_ALUctr => SEFA_ALUctr, 
--			SEFA_ExtOp => SEFA_ExtOp, 
--			SEFA_ALUSrc => SEFA_ALUSrc,
--			SEFA_MemWr => SEFA_MemWr,
--			SEFA_MemtoReg => SEFA_MemtoReg,
--			SEFA_PCSrc  => SEFA_PCSrc,
--			SEFA_RegDst => SEFA_RegDst,
--			SEFA_RegWr => SEFA_RegWr,
--);
--	
	
	GET_RegDest_Register: SEFA_SELECT_REGISTER_FILE_INPUT PORT MAP (
											SEFA_RT => SEFA_RT,
											SEFA_RD => SEFA_RD, 
											SEFA_RegDst => SEFA_RegDst,
											SEFA_REGISTER_FILE_SELECTED_INPUT => SEFA_REGISTER_FILE_SELECTED_INPUT
	);
	
	
	
	
	
	-- FOR THE FUNCTIONS THAT REQUIRE IMMEDIATE STUFF, THIS IS WHERE WE GET IT. 
	GET_EXTENDED_IMM: SEFA_IMMEDIATE_EXTENDER PORT MAP (
		SEFA_IMM16 => SEFA_IMM16,
		SEFA_ExtOp => SEFA_ExtOp,
		SEFA_EXTENDED_IMM => SEFA_EXTENDED_IMM
	
	);
	
	
	
	GET_ALU_INPUT_B:  SEFA_SELECT_SECOND_ALU_INPUT PORT MAP (
		SEFA_BUSB => SEFA_BUS_B, 
		SEFA_EXTENDED_IMM => SEFA_EXTENDED_IMM,
		SEFA_ALUsrc => SEFA_ALUsrc, 
		SEFA_INPUT_B => SEFA_INPUT_B
	);

	
	COMPUTE_ALU :  SEFA_ALU PORT MAP (
		SEFA_ALUctr => SEFA_ALUctr,
		SEFA_INPUT_A => SEFA_BUS_A, 
		SEFA_INPUT_B => SEFA_INPUT_B,
		SEFA_ALU_OUTPUT => SEFA_ALU_OUTPUT,
		SEFA_HI => SEFA_HI,
		SEFA_LO => SEFA_LO
	);
	
	
	HI_REGISTER : SEFA_HI_REGISTER PORT MAP (
		SEFA_clk => SEFA_CLOCK,
		SEFA_wren => '1',
		SEFA_rden => '1',
		SEFA_chen => '1',
		SEFA_data => SEFA_HI, 
		SEFA_HI => SEFA_HI_REGISTER_VALUE
	
	);
	
	LOW_REGISTER : SEFA_LO_REGISTER PORT MAP (
		SEFA_clk => SEFA_CLOCK,
		SEFA_wren => '1',
		SEFA_rden => '1',
		SEFA_chen => '1',
		SEFA_data => SEFA_LO, 
		SEFA_LO => SEFA_LO_REGISTER_VALUE

	);
	
	
	
	
	
	COMPUTE_DATA_MEM_COMPONET:  SEFA_NON_LPM_DATA_MEMORY PORT MAP 
	(
		SEFA_address => SEFA_ALU_OUTPUT(3 downto 0), 
		SEFA_clock => SEFA_CLOCK,
		SEFA_data => SEFA_BUS_B,
		SEFA_wren => SEFA_MemWr, 
		SEFA_q => SEFA_DATA_MEM_OUTPUT
	);
	
	COMPUTE_BUS_W_VALUE : SEFA_SELECT_MEM_TO_REG PORT MAP 
	(
		SEFA_ALU_OUTPUT => SEFA_ALU_OUTPUT,
		SEFA_DATA_MEM_OUTPUT => SEFA_DATA_MEM_OUTPUT,
		SEFA_MemtoReg => SEFA_MemtoReg, 
		SEFA_MEM_TO_REG_OUTPUT => SEFA_BUS_W
	);

	Three_Port_Ram_FINAL_RESULT : SEFA_NON_LPM_REGISTER_FILE PORT MAP (
		SEFA_clock => SEFA_CLOCK,
		SEFA_data => SEFA_BUS_W, -- TBD. what is the data supposed to be if we dont have any wtf? 
		-- isnt the purpose of this file to get it? 
		SEFA_rdaddress_a => SEFA_RS,
		SEFA_rdaddress_b => SEFA_RT,
		SEFA_wraddress => SEFA_REGISTER_FILE_SELECTED_INPUT,
		--SEFA_wren => SEFA_RegWr, 
		SEFA_wren => SEFA_RegWr, -- SHOULD BE 1 FOR LW?
		SEFA_qa => SEFA_BUS_A,
		SEFA_qb => SEFA_BUS_B
	);
	
	-- FOR BEQ AND BNE WE COMPARE R[RS] AND R[RT]
	GET_PC_COND : SEFA_Comparator_N PORT MAP ( 
			SEFA_IN0 => SEFA_BUS_A, 
			SEFA_IN1 => SEFA_BUS_B,
			SEFA_OUT => SEFA_PC_COND
	);
				
	-- UTALIZING ANL FROM BRANCHING LAB EXCEPT REPLACING OPCODE WITH PCSRC		
	NAL : SEFA_NAL PORT MAP (
		SEFA_PCSrc => SEFA_PCSrc, -- THIS IS PCSRC CONTROL SIGNAL.  
		SEFA_OPCODE => SEFA_OPCODE, -- KEEPING THIS BECAUSE TIS NEEDED FOR SELECTING IMM EXTENSION SIDE, AS WELL AS IN BRANCHING. TOO MUCH TO RECONFIGRE.
		SEFA_PC_COND => SEFA_PC_COND, -- THIS IS THE COMPARATOR CONDITION. 
		SEFA_PC_OLD => SEFA_PC,
		SEFA_IMM16 => SEFA_IMM16,
		SEFA_IMM26 => SEFA_IMM26,
		SEFA_UPDATED_PC => SEFA_PC_NEXT
	);

	
	
	

END SYN;