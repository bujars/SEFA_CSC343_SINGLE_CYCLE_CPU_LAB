LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.ALL;


ENTITY SEFA_NON_LPM_DATA_MEMORY IS
PORT(
	SEFA_clock: IN STD_LOGIC;
	SEFA_data: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	SEFA_address: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	SEFA_wren: IN STD_LOGIC;
	SEFA_q: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_NON_LPM_DATA_MEMORY;

ARCHITECTURE ARCH OF SEFA_NON_LPM_DATA_MEMORY IS
	TYPE SEFA_MEMORY IS ARRAY(0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	-- HERE WE STORE OUR VALUES IN MEMORY. NOTE THIS IS WHAT LW PULLS. THESE ARE UNIQUE AND MUST BE CHANGED TO TEST 
	-- DIFFERENT NUMBERS. 
	SIGNAL SEFA_MEM: SEFA_MEMORY := (
	 X"00000002",  
	 X"00000004",
	 X"00000006",
	 X"00000008",
	 X"0000000a",
	 X"0000000c",
	 X"0000000e",
	 X"00000010",
	 X"00000012",
	 X"00000014",
	 OTHERS => X"00000000");	
BEGIN
	PROCESS(SEFA_clock)
	 BEGIN
		IF (SEFA_clock'EVENT AND SEFA_clock = '1') THEN
			IF(SEFA_wren = '1') THEN
			SEFA_MEM(TO_INTEGER(UNSIGNED(SEFA_address))) <= SEFA_data;
		END IF;
	END IF;
	END PROCESS;
	SEFA_q <= SEFA_MEM(TO_INTEGER(UNSIGNED(SEFA_address)));
END ARCH;

