library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

-- THIS IS TO EXTEND THE IMMEDIATE FIELDS
-- BOTH SIGN AND ZERO
-- PASS INTO MUX TO DETERMINE WHICH ONE WE NEED
-- AND RETURN THE APPROPRIATE EXTENDED-IMM


-- CURRENTLY I ONLY HAVE THIS FOR IMM16 AS SEEN IN THE DIAGRAM. 

ENTITY SEFA_IMMEDIATE_EXTENDER IS
PORT(
		SEFA_IMM16 : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
		SEFA_ExtOp : IN STD_LOGIC;
		SEFA_EXTENDED_IMM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_IMMEDIATE_EXTENDER;

ARCHITECTURE ARCH OF SEFA_IMMEDIATE_EXTENDER IS
	
	SIGNAL ZERO_EXTENDED_IMM : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SIGN_EXTENDED_IMM : STD_LOGIC_VECTOR(31 DOWNTO 0);
	
BEGIN
	ZERO_EXTEND: SEFA_ZERO_EXTEND_IMM_16_TO_32 PORT MAP(
		SEFA_IMM16 => SEFA_IMM16,
		SEFA_IMM32 => ZERO_EXTENDED_IMM
	);
	
	SIGN_EXTEND: SEFA_SIGN_EXTEND_IMM_16_TO_32 PORT MAP(
		SEFA_IMM16 => SEFA_IMM16,
		SEFA_IMM32 => SIGN_EXTENDED_IMM
	);
	
	EXTEND_MUX: SEFA_IMMEDIATE_EXTENDED_MUX PORT MAP(
		SEFA_ZERO_EXTENDED_IMM => ZERO_EXTENDED_IMM,
		SEFA_SIGN_EXTENDED_IMM => SIGN_EXTENDED_IMM,
		SEFA_ExtOp => SEFA_ExtOp, 
		SEFA_EXTENDED_IMM => SEFA_EXTENDED_IMM
	
	);
	
END ARCH;
