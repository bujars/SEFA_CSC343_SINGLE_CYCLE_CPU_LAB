LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.ALL;


-- THIS IS THE FILE THAT COMPUTES AND OF INPUT A AND INPUT B


ENTITY SEFA_AND_COMPONENT IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_AND_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
);
END SEFA_AND_COMPONENT;

ARCHITECTURE ARCH OF SEFA_AND_COMPONENT IS
BEGIN
	
	SEFA_AND_RESULT <= SEFA_INPUT_A AND SEFA_INPUT_B;

END ARCH;