library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

-- THIS IS TO CHOOSE THE SECOND DATA INPUT INTO
-- ALU based on ALUsrc value
-- THIS IS A 2-1 MULTIPLEXER WHERE ALUsrc IS THE SELECT BIT


ENTITY SEFA_SELECT_SECOND_ALU_INPUT IS
PORT(
		SEFA_BUSB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_EXTENDED_IMM : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_ALUsrc : IN STD_LOGIC;
		SEFA_INPUT_B : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_SELECT_SECOND_ALU_INPUT;

ARCHITECTURE ARCH OF SEFA_SELECT_SECOND_ALU_INPUT IS
	
BEGIN


	SEFA_INPUT_B <= SEFA_EXTENDED_IMM WHEN SEFA_ALUsrc = '1' 
							ELSE SEFA_BUSB;

END ARCH;
