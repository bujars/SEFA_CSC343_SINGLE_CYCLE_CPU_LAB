library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;


-- The purpose of this component is to select between PC+4 or PC+SignExtended(Imm16)+4 OR PC+SIGNEXTENDED(IMM26)+4
-- It must call the appropriate components that perform the addtion.

-- NOTE, HERE WE HANDLE THE PC INCREMENTING LOGIC BASED ON
-- OPCODE AND RS, RT COMPARISON (FOR BEQ AND BNE)
-- OPCODE: 000100 = BEQ
-- OPCODE: 000101 = BNE
-- OPCODE: 000010 = J 

-- *OPCODES COME FROM THE MIPS GREEN PAGES: https://courses.cs.washington.edu/courses/cse378/09au/MIPS_Green_Sheet.pdf

-- NOTE, I MIGHT NEED TO REVIST BECAUSE OF THE PCSRC... CONTROL SIGNAL...(BUT MIGHT JUST BE PC SELECTOR -- NO THIS IS FOR BEQ VS BNE)

ENTITY SEFA_BRANCHING_MUX IS
	PORT(
		SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		SEFA_PC_Plus_4 : IN STD_LOGIC_VECTOR(31 DOWNTo 0);
		SEFA_PC_IMM_Plus_4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_PC_SELECTOR : IN STD_LOGIC; 
		SEFA_PC_NEW : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END SEFA_BRANCHING_MUX;

ARCHITECTURE arch OF SEFA_BRANCHING_MUX IS
BEGIN
	SEFA_PC_NEW <= SEFA_PC_IMM_Plus_4 WHEN 
									(SEFA_OPCODE = "000010"  -- J
									OR (SEFA_PC_SELECTOR = '1'   AND  SEFA_OPCODE = "000100"   ) -- BEQ
									OR (SEFA_PC_SELECTOR = '0' AND SEFA_OPCODE = "000101") -- BNE
									)
							ELSE SEFA_PC_Plus_4;

END arch;