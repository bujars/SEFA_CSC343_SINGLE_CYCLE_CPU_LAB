library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

-- THIS IS TO CHOOSE THE INPUT TO REGISTERS FILE
-- IE RT OR RD
-- BASED ON RegDst


ENTITY SEFA_SELECT_REGISTER_FILE_INPUT IS
PORT(
		SEFA_RT: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		SEFA_RD : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		SEFA_RegDst : IN STD_LOGIC;
		SEFA_REGISTER_FILE_SELECTED_INPUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
);
END SEFA_SELECT_REGISTER_FILE_INPUT;

ARCHITECTURE ARCH OF SEFA_SELECT_REGISTER_FILE_INPUT IS
	
BEGIN


	SEFA_REGISTER_FILE_SELECTED_INPUT <= SEFA_RD WHEN SEFA_RegDst = '1' 
							ELSE SEFA_RT;

END ARCH;
