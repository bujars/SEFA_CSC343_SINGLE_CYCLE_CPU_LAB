LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.ALL;


-- THIS IS THE FILE THAT CHOOSES WHICH OPERATION THE ALU IS SUPPOSED TO OUTPUT. 
-- IT TAKES IN ALL THE RESULTS OF THE DIFFERNT ALU OPERATIONS AND SELECTS THE OUTPUT USING WHEN CLAUSE WITH CODE CONDITION CHECKING.


ENTITY SEFA_ALU_MUX IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_CONDITION_CODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_ADD : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_SUB : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ALU_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
	-- NOTE IM NOT SURE HOW WE ARE GOING TO DO OUTPUT FOR MUL/DIV WHICH IS 64 BITS.......FOR NOW IGNORING.
	-- pOSSIBLY HAVE TWO OUTPUTS ONE
	-- MULT: FIRST HAS FIRST 32 BITS SECOND HAS SECOND 32 BITS
	-- DIV: FIRST HAS QUOT SECOND HAS REMAINDER
	-- FOR OTHER OPERATIONS WE ONLY FOCUS ON MAIN ONE. 
);
END SEFA_ALU_MUX;

ARCHITECTURE ARCH OF SEFA_ALU_MUX IS
BEGIN
	
	SEFA_ALU_RESULT <= SEFA_ADD WHEN SEFA_CONDITION_CODE = "000000"
							ELSE SEFA_SUB;


END ARCH;