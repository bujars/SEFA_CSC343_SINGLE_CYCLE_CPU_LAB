LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE SEFA_SINGLE_CYCLE_CPU_PACKAGE IS

COMPONENT SEFA_ALU IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_FUNCT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ALU_OUTPUT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
	-- NOTE IM NOT SURE HOW WE ARE GOING TO DO OUTPUT FOR MUL/DIV WHICH IS 64 BITS.......FOR NOW IGNORING.
);
END COMPONENT SEFA_ALU;

COMPONENT SEFA_ALU_MUX IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_FUNCT: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	SEFA_ADD : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_SUB : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ADDU : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ADDI : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ADDIU : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_SUBU : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_AND : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_OR : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_NOR : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ANDI : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ORI : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_ALU_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
	-- NOTE IM NOT SURE HOW WE ARE GOING TO DO OUTPUT FOR MUL/DIV WHICH IS 64 BITS.......FOR NOW IGNORING.
);
END COMPONENT SEFA_ALU_MUX;

COMPONENT SEFA_SIGNED_LPM_ADD_SUB IS
	PORT
	(
		SEFA_add_sub		: IN STD_LOGIC ;
		SEFA_dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_overflow		: OUT STD_LOGIC ;
		SEFA_result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_SIGNED_LPM_ADD_SUB;

COMPONENT SEFA_UNSIGNED_LPM_ADD_SUB IS
	PORT
	(
		SEFA_add_sub		: IN STD_LOGIC ;
		SEFA_dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_UNSIGNED_LPM_ADD_SUB;

COMPONENT SEFA_AND_COMPONENT IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_AND_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
);
END COMPONENT SEFA_AND_COMPONENT;

COMPONENT SEFA_OR_COMPONENT IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_OR_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
);
END COMPONENT SEFA_OR_COMPONENT;

COMPONENT SEFA_NOR_COMPONENT IS 
GENERIC(SEFA_N : INTEGER := 32);
PORT(
	SEFA_INPUT_A : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_INPUT_B : IN STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0);
	SEFA_NOR_RESULT : OUT STD_LOGIC_VECTOR(SEFA_N-1 DOWNTO 0)
);
END COMPONENT SEFA_NOR_COMPONENT;

COMPONENT SEFA_LPM_MULT IS
	PORT
	(
		SEFA_dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
END COMPONENT SEFA_LPM_MULT;

COMPONENT SEFA_LPM_DIVIDE IS
	PORT
	(
		SEFA_denom		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_numer		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_quotient		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		SEFA_remain		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END COMPONENT SEFA_LPM_DIVIDE;


COMPONENT SEFA_Register_N_VHDL is 
	generic (SEFA_N: integer := 32); -- The genetics feature permits us to change the side of this register desin easily. Its a const variable
	port (
		SEFA_clk: in std_logic; -- clock
		SEFA_wren: in std_logic; -- write enable (if it is 0, the stored data will not change)
		SEFA_rden: in std_logic; -- read enable (only when it is 1, the stored data will be displayed to output)
		SEFA_chen: in std_logic; --  chip enable (if it is 0, the output will be undefined)
		SEFA_data: in std_logic_vector (SEFA_N-1 downto 0); -- data input
		SEFA_q: out std_logic_vector(SEFA_N-1 downto 0) -- output. This is essentially just a display
		);
end COMPONENT SEFA_Register_N_VHDL;


COMPONENT SEFA_IR_REGISTER IS
	generic (SEFA_N: integer := 32);
	port(
	SEFA_clk: in std_logic; -- clock
		SEFA_wren: in std_logic; -- write enable (if it is 0, the stored data will not change)
		SEFA_rden: in std_logic; -- read enable (only when it is 1, the stored data will be displayed to output)
		SEFA_chen: in std_logic; --  chip enable (if it is 0, the output will be undefined)
		SEFA_data: in std_logic_vector (SEFA_N-1 downto 0); -- data input
		SEFA_IR: out std_logic_vector(SEFA_N-1 downto 0)
		);
end COMPONENT SEFA_IR_REGISTER;



END SEFA_SINGLE_CYCLE_CPU_PACKAGE;