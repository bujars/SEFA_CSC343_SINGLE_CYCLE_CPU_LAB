library IEEE;
use IEEE.std_logic_1164.all;
use work.SEFA_SINGLE_CYCLE_CPU_PACKAGE.all;

-- THIS IS TO CHOOSE THE DATA that goes back to the registers after we finish ALU + Data Mem
-- We select based on MemtoReg control signal. 

ENTITY SEFA_SELECT_MEM_TO_REG IS
PORT(
		SEFA_ALU_OUTPUT: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_DATA_MEM_OUTPUT : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEFA_MemtoReg : IN STD_LOGIC;
		SEFA_MEM_TO_REG_OUTPUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END SEFA_SELECT_MEM_TO_REG;

ARCHITECTURE ARCH OF SEFA_SELECT_MEM_TO_REG IS
	
BEGIN


	SEFA_MEM_TO_REG_OUTPUT <= SEFA_DATA_MEM_OUTPUT WHEN SEFA_MemtoReg = '1' 
							ELSE SEFA_ALU_OUTPUT;

END ARCH;
